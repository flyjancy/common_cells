// -----------------------------Details----------------------------------- // 
// File        : uart_tx.v
// Author      : pastglory
// Date        : 
// Version     : 1.0
// Description : transfor data
// -----------------------------History----------------------------------- //
// Date      BY          Version  Change Description
//
//   pastglory   1.0      Initial Release. 
// ----------------------------------------------------------------------- // 

module uart_tx (
    //TODO
);

endmodule