// -----------------------------Details----------------------------------- // 
// File        : uart_tx.v
// Author      : pastglory
// Date        : 
// Version     : 1.0
// Description : transfor data
// -----------------------------History----------------------------------- //
// Date      BY          Version  Change Description
//
//   pastglory   1.0      Initial Release. 
// ----------------------------------------------------------------------- // 

module uart_tx (
    input           clk,        // fpga clock
    input           clk_uart,   // UART clock
    input           rst_n,      // reset
    input [7 : 0]   data,       // data for trans
    output          txd         // tx data
);

//TODO

endmodule